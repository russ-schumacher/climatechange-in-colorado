netcdf tmp_mask.baseflow {
dimensions:
	Lon = 12 ;
	Lat = 16 ;
	Time = UNLIMITED ; // (1 currently)
variables:
	float Lon(Lon) ;
		Lon:long_name = "longitude" ;
		Lon:standard_name = "longitude" ;
		Lon:units = "degreesE" ;
	float Lat(Lat) ;
		Lat:long_name = "latitude" ;
		Lat:standard_name = "latitude" ;
		Lat:units = "degreesN" ;
	double Time(Time) ;
		Time:long_name = "time" ;
		Time:units = "days since 1800-01-01" ;
	float baseflow(Time, Lat, Lon) ;
		baseflow:long_name = "baseflow" ;
		baseflow:units = "mm/day" ;
		baseflow:missing_value = 1.e+30f ;
		baseflow:_FillValue = 1.e+30f ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:creation_date = "Fri Jul 15 12:45:58 2016" ;
		:output_version = 0 ;
		:version_description = "" ;
		:created_by = "pierce" ;
		:cmd_line = "/home/pierce/src/mine/vic_utils/xtslab2nc -rm_slabs -template /net/loca2/LOCA_2016-04-02/ACCESS1-0/16th/historical/r1i1p1/tasmax/tasmax_day_ACCESS1-0_historical_r1i1p1_20050101-20051231.LOCA_2016-04-02.16th.nc -dir ../vic_output.historical -fname_base flux_snow -flux ../../fluxdescrip_dpierce_27_vars.txt" ;
		:run_in_directory = "/home/pierce/projects/vic_LOCA/NAmer/ACCESS1-0/vic_output.historical.netcdf" ;
data:

 Lon = -106.5938, -106.5312, -106.4688, -106.4062, -106.3438, -106.2812, 
    -106.2188, -106.1562, -106.0938, -106.0312, -105.9688, -105.9062 ;

 Lat = 38.40625, 38.46875, 38.53125, 38.59375, 38.65625, 38.71875, 38.78125, 
    38.84375, 38.90625, 38.96875, 39.03125, 39.09375, 39.15625, 39.21875, 
    39.28125, 39.34375 ;

 Time = 54786 ;

 baseflow =
   _, _, _, _, _, _, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, 1, 1, 1, 1, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, 
   1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, _, _, _, _ ;
}
