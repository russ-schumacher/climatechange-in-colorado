netcdf tmp_mask.SWE {
dimensions:
	Lon = 24 ;
	Lat = 18 ;
	Time = UNLIMITED ; // (1 currently)
variables:
	float Lon(Lon) ;
		Lon:long_name = "longitude" ;
		Lon:standard_name = "longitude" ;
		Lon:units = "degreesE" ;
	float Lat(Lat) ;
		Lat:long_name = "latitude" ;
		Lat:standard_name = "latitude" ;
		Lat:units = "degreesN" ;
	double Time(Time) ;
		Time:long_name = "time" ;
		Time:units = "days since 1800-01-01" ;
	float SWE(Time, Lat, Lon) ;
		SWE:long_name = "snow_water_equivalent" ;
		SWE:units = "mm" ;
		SWE:missing_value = 1.e+30f ;
		SWE:_FillValue = 1.e+30f ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:creation_date = "Fri Jul 15 14:30:43 2016" ;
		:output_version = 0 ;
		:version_description = "" ;
		:created_by = "pierce" ;
		:cmd_line = "/home/pierce/src/mine/vic_utils/xtslab2nc -rm_slabs -template /net/loca2/LOCA_2016-04-02/ACCESS1-0/16th/historical/r1i1p1/tasmax/tasmax_day_ACCESS1-0_historical_r1i1p1_20050101-20051231.LOCA_2016-04-02.16th.nc -dir ../vic_output.historical -fname_base flux_snow -flux ../../fluxdescrip_dpierce_27_vars.txt" ;
		:run_in_directory = "/home/pierce/projects/vic_LOCA/NAmer/ACCESS1-0/vic_output.historical.netcdf" ;
data:

 Lon = -107.7188, -107.6562, -107.5938, -107.5312, -107.4688, -107.4062, 
    -107.3438, -107.2812, -107.2188, -107.1562, -107.0938, -107.0312, 
    -106.9688, -106.9062, -106.8438, -106.7812, -106.7188, -106.6562, 
    -106.5938, -106.5312, -106.4688, -106.4062, -106.3438, -106.2812 ;

 Lat = 37.90625, 37.96875, 38.03125, 38.09375, 38.15625, 38.21875, 38.28125, 
    38.34375, 38.40625, 38.46875, 38.53125, 38.59375, 38.65625, 38.71875, 
    38.78125, 38.84375, 38.90625, 38.96875 ;

 Time = 54786 ;

 SWE =
   _, _, _, _, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, 
   _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
   _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, 
   _, _, _, _, _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _ ;
}
