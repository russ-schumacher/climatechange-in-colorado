netcdf tmp_mask.baseflow {
dimensions:
	Lon = 18 ;
	Lat = 10 ;
	Time = UNLIMITED ; // (1 currently)
variables:
	float Lon(Lon) ;
		Lon:long_name = "longitude" ;
		Lon:standard_name = "longitude" ;
		Lon:units = "degreesE" ;
	float Lat(Lat) ;
		Lat:long_name = "latitude" ;
		Lat:standard_name = "latitude" ;
		Lat:units = "degreesN" ;
	double Time(Time) ;
		Time:long_name = "time" ;
		Time:units = "days since 1800-01-01" ;
	float baseflow(Time, Lat, Lon) ;
		baseflow:long_name = "baseflow" ;
		baseflow:units = "mm/day" ;
		baseflow:missing_value = 1.e+30f ;
		baseflow:_FillValue = 1.e+30f ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:creation_date = "Fri Jul 15 12:45:58 2016" ;
		:output_version = 0 ;
		:version_description = "" ;
		:created_by = "pierce" ;
		:cmd_line = "/home/pierce/src/mine/vic_utils/xtslab2nc -rm_slabs -template /net/loca2/LOCA_2016-04-02/ACCESS1-0/16th/historical/r1i1p1/tasmax/tasmax_day_ACCESS1-0_historical_r1i1p1_20050101-20051231.LOCA_2016-04-02.16th.nc -dir ../vic_output.historical -fname_base flux_snow -flux ../../fluxdescrip_dpierce_27_vars.txt" ;
		:run_in_directory = "/home/pierce/projects/vic_LOCA/NAmer/ACCESS1-0/vic_output.historical.netcdf" ;
data:

 Lon = -107.4688, -107.4062, -107.3438, -107.2812, -107.2188, -107.1562, 
    -107.0938, -107.0312, -106.9688, -106.9062, -106.8438, -106.7812, 
    -106.7188, -106.6562, -106.5938, -106.5312, -106.4688, -106.4062 ;

 Lat = 37.40625, 37.46875, 37.53125, 37.59375, 37.65625, 37.71875, 37.78125, 
    37.84375, 37.90625, 37.96875 ;

 Time = 54786 ;

 baseflow =
   _, _, _, _, _, _, _, _, _, _, _, _, 1, 1, _, _, _, _, 
   _, _, _, _, _, _, _, _, _, _, _, _, 1, 1, _, _, _, _, 
   _, _, _, _, _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 
   _, _, _, _, _, _, _, _, _, _, 1, 1, 1, 1, 1, 1, 1, 1, 
   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, _, _, 
   _, _, _, _, _, _, 1, 1, 1, 1, _, _, _, _, _, _, _, _, 
   _, _, _, _, _, _, 1, 1, 1, 1, _, _, _, _, _, _, _, _ ;
}
